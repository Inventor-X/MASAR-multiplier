`timescale 1ns / 1ps

module masar_tb(

    );
    reg [7:0] x,y;
    wire[15:0] result;

    
    //temperory outputs 
    masar DUT(x,y,result);
    initial begin
        x<= 16'd55;
        y<= 16'd63;
    #30 x<=16'd22;
        y<=16'd3;
    #30 x<=16'd23;
        y<=16'd69;
    #30 x<=16'd55;
        y<=16'd62;
    #30 x<=16'd12;
        y<=16'd34;
    #30 x<=16'd126;
        y<=16'd69;
    #30 x<=16'd28;
        y<=16'd32;
    #30 x<=16'd60;
        y<=16'd24;
    #30 x<=16'd48;
        y<=16'd12;
    #30 x<=16'd482;
        y<=16'd124;
    #30 x<=16'd485;
        y<=16'd127;
    #30 x<=16'd23;
        y<=16'd124;
    #30 x<=16'd485;
        y<=16'd122;
    #30 x<=16'd126;
        y<=16'd125;
    #30 x<= 16'd55;
        y<= 16'd789;
    #30 x<=16'd233;
        y<=16'd64;
    #30 x<=16'd53;
        y<=16'd89;
    #30 x<=16'd15;
        y<=16'd452;
    #30 x<=16'd122;
        y<=16'd343;
    #30 x<=16'd126;
        y<=16'd693;
    #30 x<=16'd280;
        y<=16'd324;
    #30 x<=16'd600;
        y<=16'd243;
    #30 x<=16'd480;
        y<=16'd121;
    #30 x<=16'd482;
        y<=16'd124;
    #30 x<=16'd485;
        y<=16'd127;
    #30 x<=16'd23;
        y<=16'd124;
    #30 x<=16'd485;
        y<=16'd122;
    #30 x<=16'd126;
        y<=16'd125;
    #30 x<=16'd0;
        y<=16'd0;
        
       
    end
    
endmodule
